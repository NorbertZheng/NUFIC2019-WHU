`timescale 1ns/1ns
module test_ThresholdCutter #(
	parameter		// config enable
					CONFIG_EN							=	0,		// do not enable config
					// config
					CLK_FRE								=	50,		// 50MHz
					BAUD_RATE							=	115200,	// 115200Hz (4800, 19200, 38400, 57600, 115200, 38400...)
					STOP_BIT							=	0,		// 0 : 1-bit stop-bit, 1 : 2-bit stop-bit
					CHECK_BIT							=	0,		// 0 : no check-bit, 1 : odd, 2 : even
					// default	9600	0	0
					// granularity
					REQUEST_FIFO_DATA_WIDTH				=	8,		// the bit width of data we stored in the FIFO
					REQUEST_FIFO_DATA_DEPTH_INDEX		=	5,		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
					RESPONSE_FIFO_DATA_WIDTH			=	8,		// the bit width of data we stored in the FIFO
					RESPONSE_FIFO_DATA_DEPTH_INDEX		=	5,		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
					// uart connected with PC
					PC_BAUD_RATE						=	115200,	// 115200Hz
					// enable simulation
					SIM_ENABLE							=	1,				// enable simulation
					// parameter for window
					WINDOW_DEPTH_INDEX					=	7,				// support up to 128 windows
					WINDOW_DEPTH						=	100,			// 100 windows
					WINDOW_WIDTH						=	(32 << 3),		// 32B window
					THRESHOLD							=	32'h0010_0000,	// threshold
					BLOCK_NUM_INDEX						=	4,				// 2 ** 6 == 64 blocks		// 16
					// parameter for package
					A_OFFSET							=	2,				// A's offset
					// parameter for square
					SQUARE_SRC_DATA_WIDTH				=	16,				// square src data width
					// parameter for preset-sequence
					PRESET_SEQUENCE						=	128'h00_01_02_03_04_05_06_07_08_09_00_01_02_03_04_05,
					// parameter for package
					PACKAGE_SIZE						=	11,
					PACKAGE_NUM							=	4,
					// parameter for uart
					TX_DATA_BYTE_WIDTH					=	11,		// 11 bytes to transmit
					RX_DATA_BYTE_WIDTH					=	11		// 11 bytes to receive
	`ifndef			TX_DATA_BIT_WIDTH
	`define			TX_DATA_BIT_WIDTH					(TX_DATA_BYTE_WIDTH << 3)
	`endif
	`ifndef			RX_DATA_BIT_WIDTH
	`define			RX_DATA_BIT_WIDTH					(RX_DATA_BYTE_WIDTH << 3)
	`endif
) (

);

	reg clk, rst_n;
	// ThresholdCutter signals
	wire BlueTooth_Txd;
	// sim_BlueTooth signals
	wire uart_tx;
	reg tx_vld;
	reg [`TX_DATA_BIT_WIDTH - 1:0] tx_data;

	// testsuite
	always # 50
		clk = ~clk;

	initial
		begin
		clk = 1'b0;
		rst_n = 1'b1;
		tx_vld = 1'b0;
		tx_data = {WINDOW_WIDTH{1'b0}};
		# 500;
		rst_n = 1'b0;
		# 500;
		rst_n = 1'b1;
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 39900;		// 400 - period
		end

	// sim_BlueTooth
	sim_BlueTooth #(
		// config
		.CLK_FRE(CLK_FRE),		// 50MHz
		.BAUD_RATE(BAUD_RATE),	// 9600Hz (4800, 19200, 38400, 57600, 115200, 38400...)
		.TX_DATA_BYTE_WIDTH(TX_DATA_BYTE_WIDTH),	// 11 bytes to transmit
		.RX_DATA_BYTE_WIDTH(RX_DATA_BYTE_WIDTH)		// 11 bytes to receive
	) m_sim_BlueTooth (
		.clk				(clk			),
		.rst_n				(rst_n			),

		// uart signals
		.uart_rx			(				),
		.uart_tx			(uart_tx		),		// should connect with BlueTooth_Txd in BlueToothController.v

		// inner data
		.tx_data			(tx_data		),		// data
		.tx_vld				(tx_vld			),		// start the transmit process
		.tx_rdy				(				),		// transmit process complete
		.rx_data			(				),		// data
		.rx_ack				(				),		// data is received by receiver buffer					(RX_WAIT)
		.rx_rdy				(				)		// send signal to receiver buffer that data is ready
	);

	// ThresholdCutter
	ThresholdCutter #(
		// config enable
		.CONFIG_EN(CONFIG_EN),		// do not enable config
		// config
		.CLK_FRE(CLK_FRE),		// 50MHz
		.BAUD_RATE(BAUD_RATE),	// 115200Hz (4800, 19200, 38400, 57600, 115200, 38400...)
		.STOP_BIT(STOP_BIT),		// 0 : 1-bit stop-bit, 1 : 2-bit stop-bit
		.CHECK_BIT(CHECK_BIT),		// 0 : no check-bit, 1 : odd, 2 : even
		// default	9600	0	0
		// granularity
		.REQUEST_FIFO_DATA_WIDTH(REQUEST_FIFO_DATA_WIDTH),		// the bit width of data we stored in the FIFO
		.REQUEST_FIFO_DATA_DEPTH_INDEX(REQUEST_FIFO_DATA_DEPTH_INDEX),		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
		.RESPONSE_FIFO_DATA_WIDTH(RESPONSE_FIFO_DATA_WIDTH),		// the bit width of data we stored in the FIFO
		.RESPONSE_FIFO_DATA_DEPTH_INDEX(RESPONSE_FIFO_DATA_DEPTH_INDEX),		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
		// uart connected with PC
		.PC_BAUD_RATE(PC_BAUD_RATE),	// 115200Hz
		// enable simulation
		.SIM_ENABLE(SIM_ENABLE),				// enable simulation
		// parameter for window
		.WINDOW_DEPTH_INDEX(WINDOW_DEPTH_INDEX),				// support up to 128 windows
		.WINDOW_DEPTH(WINDOW_DEPTH),			// 100 windows
		.WINDOW_WIDTH(WINDOW_WIDTH),		// 32B window
		.THRESHOLD(THRESHOLD),	// threshold
		.BLOCK_NUM_INDEX(BLOCK_NUM_INDEX),				// 2 ** 6 == 64 blocks		// 16
		// parameter for package
		.A_OFFSET(A_OFFSET),				// A's offset
		// parameter for square
		.SQUARE_SRC_DATA_WIDTH(SQUARE_SRC_DATA_WIDTH),				// square src data width
		// parameter for preset-sequence
		.PRESET_SEQUENCE(PRESET_SEQUENCE),
		// parameter for package
		.PACKAGE_SIZE(PACKAGE_SIZE),
		.PACKAGE_NUM(PACKAGE_NUM)
	) m_ThresholdCutter (
		.clk							(clk				),
		.rst_n							(rst_n				),

		// BlueTooth_Config
		.BlueTooth_State				(					),
		.BlueTooth_Key					(					),
		.BlueTooth_Rxd					(					),
		.BlueTooth_Txd					(BlueTooth_Txd		),
		.BlueTooth_Vcc					(					),
		.BlueTooth_Gnd					(					),

		// ThresholdCutterWindow signals
		.ThresholdCutterWindow_flag_o	(					),

		// AXI RAM signals
		// ram safe access
		.rsta_busy						(					),
		.rstb_busy						(					),

		// AXI read control signals
		.s_axi_arid						(					),
		.s_axi_araddr					(					),
		.s_axi_arlen					(					),
		.s_axi_arsize					(					),
		.s_axi_arburst					(					),
		.s_axi_arvalid					(					),
		.s_axi_arready					(					),

		// AXI read data signals
		.s_axi_rid						(					),
		.s_axi_rdata					(					),
		.s_axi_rresp					(					),
		.s_axi_rlast					(					),
		.s_axi_rvalid					(					),
		.s_axi_rready					(					)
	);
	assign BlueTooth_Txd = uart_tx;

endmodule
