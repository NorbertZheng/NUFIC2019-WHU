`timescale 1ns/1ns
module test_ThresholdCutterWindow #(
	parameter		// enable simulation
					SIM_ENABLE				=	0,				// enable simulation
					// parameter for window
					WINDOW_DEPTH_INDEX		=	7,				// support up to 128 windows
					WINDOW_DEPTH			=	100,			// 100 windows
					WINDOW_WIDTH			=	(32 << 3),		// 32-B window
					THRESHOLD				=	32'h0010_0000,	// threshold
					BLOCK_NUM_INDEX			=	4,				// 2 ** 6 == 64 blocks
					// parameter for package
					A_OFFSET				=	2,				// A's offset
					// parameter for square
					SQUARE_SRC_DATA_WIDTH	=	16,				// square src data width
					// parameter for preset-sequence
					PRESET_SEQUENCE			=	128'h00_01_02_03_04_05_06_07_08_09_00_01_02_03_04_05
	`define			sim_window
) (

);

	// ThresholdCutterWindow signals
	reg clk, rst_n, data_wen;
	reg [WINDOW_WIDTH:0] data_i;
	wire [WINDOW_DEPTH - 1:0] flag_o;

	// testsuite
	always # 50
		clk = ~clk;

	initial
		begin
		clk = 1'b0;
		rst_n = 1'b1;
		data_wen = 1'b0;
		data_i = {(WINDOW_WIDTH + 1){1'b0}};
		# 500;
		rst_n = 1'b0;
		# 500;
		rst_n = 1'b1;
				data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_20_00_20_00_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_01_20_01_20_01_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_02_20_02_20_02_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_03_20_03_20_03_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_04_20_04_20_04_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_05_20_05_20_05_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_06_20_06_20_06_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_07_20_07_20_07_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_08_20_08_20_08_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_09_20_09_20_09_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0a_20_0a_20_0a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0b_20_0b_20_0b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0c_20_0c_20_0c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0d_20_0d_20_0d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0e_20_0e_20_0e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0f_20_0f_20_0f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_10_20_10_20_10_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_11_20_11_20_11_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_12_20_12_20_12_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_13_20_13_20_13_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_14_20_14_20_14_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_15_20_15_20_15_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_16_20_16_20_16_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_17_20_17_20_17_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_18_20_18_20_18_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_19_20_19_20_19_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1a_20_1a_20_1a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1b_20_1b_20_1b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1c_20_1c_20_1c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1d_20_1d_20_1d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1e_20_1e_20_1e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1f_20_1f_20_1f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_20_20_20_20_20_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_21_20_21_20_21_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_22_20_22_20_22_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_23_20_23_20_23_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_24_20_24_20_24_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_25_20_25_20_25_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_26_20_26_20_26_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_27_20_27_20_27_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_28_20_28_20_28_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_29_20_29_20_29_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2a_20_2a_20_2a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2b_20_2b_20_2b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2c_20_2c_20_2c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2d_20_2d_20_2d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2e_20_2e_20_2e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2f_20_2f_20_2f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_30_20_30_20_30_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_31_20_31_20_31_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_32_20_32_20_32_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_33_20_33_20_33_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_34_20_34_20_34_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_35_20_35_20_35_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_36_20_36_20_36_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_37_20_37_20_37_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_38_20_38_20_38_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_39_20_39_20_39_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3a_20_3a_20_3a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3b_20_3b_20_3b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3c_20_3c_20_3c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3d_20_3d_20_3d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3e_20_3e_20_3e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3f_20_3f_20_3f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_40_20_40_20_40_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_41_20_41_20_41_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_42_20_42_20_42_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_43_20_43_20_43_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_44_20_44_20_44_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_45_20_45_20_45_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_46_20_46_20_46_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_47_20_47_20_47_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_48_20_48_20_48_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_49_20_49_20_49_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4a_20_4a_20_4a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4b_20_4b_20_4b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4c_20_4c_20_4c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4d_20_4d_20_4d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4e_20_4e_20_4e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4f_20_4f_20_4f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_50_20_50_20_50_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_51_20_51_20_51_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_52_20_52_20_52_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_53_20_53_20_53_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_54_20_54_20_54_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_55_20_55_20_55_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_56_20_56_20_56_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_57_20_57_20_57_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_58_20_58_20_58_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_59_20_59_20_59_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5a_20_5a_20_5a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5b_20_5b_20_5b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5c_20_5c_20_5c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5d_20_5d_20_5d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5e_20_5e_20_5e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5f_20_5f_20_5f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_60_20_60_20_60_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_61_20_61_20_61_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_62_20_62_20_62_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_63_20_63_20_63_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_64_20_64_20_64_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_65_20_65_20_65_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_66_20_66_20_66_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_67_20_67_20_67_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_68_20_68_20_68_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_69_20_69_20_69_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6a_20_6a_20_6a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6b_20_6b_20_6b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6c_20_6c_20_6c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6d_20_6d_20_6d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6e_20_6e_20_6e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6f_20_6f_20_6f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_70_20_70_20_70_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_71_20_71_20_71_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_72_20_72_20_72_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_73_20_73_20_73_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_74_20_74_20_74_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_75_20_75_20_75_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_76_20_76_20_76_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_77_20_77_20_77_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_78_20_78_20_78_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_79_20_79_20_79_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7a_20_7a_20_7a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7b_20_7b_20_7b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7c_20_7c_20_7c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7d_20_7d_20_7d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7e_20_7e_20_7e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7f_20_7f_20_7f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_80_20_80_20_80_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_81_20_81_20_81_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_82_20_82_20_82_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_83_20_83_20_83_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_84_20_84_20_84_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_85_20_85_20_85_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_86_20_86_20_86_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_87_20_87_20_87_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_88_20_88_20_88_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_89_20_89_20_89_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8a_20_8a_20_8a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8b_20_8b_20_8b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8c_20_8c_20_8c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8d_20_8d_20_8d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8e_20_8e_20_8e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8f_20_8f_20_8f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_90_20_90_20_90_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_91_20_91_20_91_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_92_20_92_20_92_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_93_20_93_20_93_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_94_20_94_20_94_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_95_20_95_20_95_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_96_20_96_20_96_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_97_20_97_20_97_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_98_20_98_20_98_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_99_20_99_20_99_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9a_20_9a_20_9a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9b_20_9b_20_9b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9c_20_9c_20_9c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9d_20_9d_20_9d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9e_20_9e_20_9e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9f_20_9f_20_9f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a0_20_a0_20_a0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a1_20_a1_20_a1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a2_20_a2_20_a2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a3_20_a3_20_a3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a4_20_a4_20_a4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a5_20_a5_20_a5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a6_20_a6_20_a6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a7_20_a7_20_a7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a8_20_a8_20_a8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a9_20_a9_20_a9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_aa_20_aa_20_aa_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ab_20_ab_20_ab_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ac_20_ac_20_ac_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ad_20_ad_20_ad_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ae_20_ae_20_ae_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_af_20_af_20_af_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b0_20_b0_20_b0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b1_20_b1_20_b1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b2_20_b2_20_b2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b3_20_b3_20_b3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b4_20_b4_20_b4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b5_20_b5_20_b5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b6_20_b6_20_b6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b7_20_b7_20_b7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b8_20_b8_20_b8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b9_20_b9_20_b9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ba_20_ba_20_ba_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bb_20_bb_20_bb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bc_20_bc_20_bc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bd_20_bd_20_bd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_be_20_be_20_be_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bf_20_bf_20_bf_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c0_20_c0_20_c0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c1_20_c1_20_c1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c2_20_c2_20_c2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c3_20_c3_20_c3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c4_20_c4_20_c4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c5_20_c5_20_c5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c6_20_c6_20_c6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c7_20_c7_20_c7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c8_20_c8_20_c8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c9_20_c9_20_c9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ca_20_ca_20_ca_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cb_20_cb_20_cb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cc_20_cc_20_cc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cd_20_cd_20_cd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ce_20_ce_20_ce_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cf_20_cf_20_cf_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d0_20_d0_20_d0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d1_20_d1_20_d1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d2_20_d2_20_d2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d3_20_d3_20_d3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d4_20_d4_20_d4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d5_20_d5_20_d5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d6_20_d6_20_d6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d7_20_d7_20_d7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d8_20_d8_20_d8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d9_20_d9_20_d9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_da_20_da_20_da_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_db_20_db_20_db_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_dc_20_dc_20_dc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_dd_20_dd_20_dd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_de_20_de_20_de_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_df_20_df_20_df_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e0_20_e0_20_e0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e1_20_e1_20_e1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e2_20_e2_20_e2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e3_20_e3_20_e3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e4_20_e4_20_e4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e5_20_e5_20_e5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e6_20_e6_20_e6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e7_20_e7_20_e7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e8_20_e8_20_e8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e9_20_e9_20_e9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ea_20_ea_20_ea_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_eb_20_eb_20_eb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ec_20_ec_20_ec_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ed_20_ed_20_ed_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ee_20_ee_20_ee_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ef_20_ef_20_ef_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f0_20_f0_20_f0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f1_20_f1_20_f1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f2_20_f2_20_f2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f3_20_f3_20_f3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f4_20_f4_20_f4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f5_20_f5_20_f5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f6_20_f6_20_f6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f7_20_f7_20_f7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f8_20_f8_20_f8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f9_20_f9_20_f9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fa_20_fa_20_fa_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fb_20_fb_20_fb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fc_20_fc_20_fc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fd_20_fd_20_fd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fe_20_fe_20_fe_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ff_20_ff_20_ff_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b0};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_00_20_00_20_00_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_01_20_01_20_01_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_02_20_02_20_02_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_03_20_03_20_03_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_04_20_04_20_04_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_05_20_05_20_05_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_06_20_06_20_06_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_07_20_07_20_07_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_08_20_08_20_08_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_09_20_09_20_09_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0a_20_0a_20_0a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0b_20_0b_20_0b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0c_20_0c_20_0c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0d_20_0d_20_0d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0e_20_0e_20_0e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_0f_20_0f_20_0f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_10_20_10_20_10_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_11_20_11_20_11_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_12_20_12_20_12_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_13_20_13_20_13_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_14_20_14_20_14_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_15_20_15_20_15_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_16_20_16_20_16_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_17_20_17_20_17_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_18_20_18_20_18_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_19_20_19_20_19_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1a_20_1a_20_1a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1b_20_1b_20_1b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1c_20_1c_20_1c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1d_20_1d_20_1d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1e_20_1e_20_1e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_1f_20_1f_20_1f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_20_20_20_20_20_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_21_20_21_20_21_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_22_20_22_20_22_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_23_20_23_20_23_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_24_20_24_20_24_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_25_20_25_20_25_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_26_20_26_20_26_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_27_20_27_20_27_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_28_20_28_20_28_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_29_20_29_20_29_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2a_20_2a_20_2a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2b_20_2b_20_2b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2c_20_2c_20_2c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2d_20_2d_20_2d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2e_20_2e_20_2e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_2f_20_2f_20_2f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_30_20_30_20_30_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_31_20_31_20_31_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_32_20_32_20_32_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_33_20_33_20_33_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_34_20_34_20_34_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_35_20_35_20_35_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_36_20_36_20_36_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_37_20_37_20_37_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_38_20_38_20_38_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_39_20_39_20_39_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3a_20_3a_20_3a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3b_20_3b_20_3b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3c_20_3c_20_3c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3d_20_3d_20_3d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3e_20_3e_20_3e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_3f_20_3f_20_3f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_40_20_40_20_40_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_41_20_41_20_41_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_42_20_42_20_42_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_43_20_43_20_43_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_44_20_44_20_44_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_45_20_45_20_45_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_46_20_46_20_46_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_47_20_47_20_47_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_48_20_48_20_48_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_49_20_49_20_49_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4a_20_4a_20_4a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4b_20_4b_20_4b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4c_20_4c_20_4c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4d_20_4d_20_4d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4e_20_4e_20_4e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_4f_20_4f_20_4f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_50_20_50_20_50_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_51_20_51_20_51_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_52_20_52_20_52_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_53_20_53_20_53_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_54_20_54_20_54_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_55_20_55_20_55_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_56_20_56_20_56_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_57_20_57_20_57_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_58_20_58_20_58_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_59_20_59_20_59_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5a_20_5a_20_5a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5b_20_5b_20_5b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5c_20_5c_20_5c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5d_20_5d_20_5d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5e_20_5e_20_5e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_5f_20_5f_20_5f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_60_20_60_20_60_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_61_20_61_20_61_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_62_20_62_20_62_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_63_20_63_20_63_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_64_20_64_20_64_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_65_20_65_20_65_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_66_20_66_20_66_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_67_20_67_20_67_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_68_20_68_20_68_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_69_20_69_20_69_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6a_20_6a_20_6a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6b_20_6b_20_6b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6c_20_6c_20_6c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6d_20_6d_20_6d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6e_20_6e_20_6e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_6f_20_6f_20_6f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_70_20_70_20_70_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_71_20_71_20_71_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_72_20_72_20_72_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_73_20_73_20_73_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_74_20_74_20_74_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_75_20_75_20_75_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_76_20_76_20_76_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_77_20_77_20_77_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_78_20_78_20_78_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_79_20_79_20_79_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7a_20_7a_20_7a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7b_20_7b_20_7b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7c_20_7c_20_7c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7d_20_7d_20_7d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7e_20_7e_20_7e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_7f_20_7f_20_7f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_80_20_80_20_80_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_81_20_81_20_81_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_82_20_82_20_82_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_83_20_83_20_83_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_84_20_84_20_84_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_85_20_85_20_85_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_86_20_86_20_86_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_87_20_87_20_87_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_88_20_88_20_88_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_89_20_89_20_89_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8a_20_8a_20_8a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8b_20_8b_20_8b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8c_20_8c_20_8c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8d_20_8d_20_8d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8e_20_8e_20_8e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_8f_20_8f_20_8f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_90_20_90_20_90_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_91_20_91_20_91_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_92_20_92_20_92_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_93_20_93_20_93_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_94_20_94_20_94_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_95_20_95_20_95_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_96_20_96_20_96_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_97_20_97_20_97_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_98_20_98_20_98_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_99_20_99_20_99_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9a_20_9a_20_9a_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9b_20_9b_20_9b_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9c_20_9c_20_9c_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9d_20_9d_20_9d_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9e_20_9e_20_9e_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_9f_20_9f_20_9f_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a0_20_a0_20_a0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a1_20_a1_20_a1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a2_20_a2_20_a2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a3_20_a3_20_a3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a4_20_a4_20_a4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a5_20_a5_20_a5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a6_20_a6_20_a6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a7_20_a7_20_a7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a8_20_a8_20_a8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_a9_20_a9_20_a9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_aa_20_aa_20_aa_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ab_20_ab_20_ab_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ac_20_ac_20_ac_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ad_20_ad_20_ad_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ae_20_ae_20_ae_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_af_20_af_20_af_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b0_20_b0_20_b0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b1_20_b1_20_b1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b2_20_b2_20_b2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b3_20_b3_20_b3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b4_20_b4_20_b4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b5_20_b5_20_b5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b6_20_b6_20_b6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b7_20_b7_20_b7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b8_20_b8_20_b8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_b9_20_b9_20_b9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ba_20_ba_20_ba_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bb_20_bb_20_bb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bc_20_bc_20_bc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bd_20_bd_20_bd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_be_20_be_20_be_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_bf_20_bf_20_bf_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c0_20_c0_20_c0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c1_20_c1_20_c1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c2_20_c2_20_c2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c3_20_c3_20_c3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c4_20_c4_20_c4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c5_20_c5_20_c5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c6_20_c6_20_c6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c7_20_c7_20_c7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c8_20_c8_20_c8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_c9_20_c9_20_c9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ca_20_ca_20_ca_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cb_20_cb_20_cb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cc_20_cc_20_cc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cd_20_cd_20_cd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ce_20_ce_20_ce_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_cf_20_cf_20_cf_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d0_20_d0_20_d0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d1_20_d1_20_d1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d2_20_d2_20_d2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d3_20_d3_20_d3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d4_20_d4_20_d4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d5_20_d5_20_d5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d6_20_d6_20_d6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d7_20_d7_20_d7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d8_20_d8_20_d8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_d9_20_d9_20_d9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_da_20_da_20_da_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_db_20_db_20_db_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_dc_20_dc_20_dc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_dd_20_dd_20_dd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_de_20_de_20_de_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_df_20_df_20_df_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e0_20_e0_20_e0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e1_20_e1_20_e1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e2_20_e2_20_e2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e3_20_e3_20_e3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e4_20_e4_20_e4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e5_20_e5_20_e5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e6_20_e6_20_e6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e7_20_e7_20_e7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e8_20_e8_20_e8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_e9_20_e9_20_e9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ea_20_ea_20_ea_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_eb_20_eb_20_eb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ec_20_ec_20_ec_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ed_20_ed_20_ed_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ee_20_ee_20_ee_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ef_20_ef_20_ef_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f0_20_f0_20_f0_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f1_20_f1_20_f1_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f2_20_f2_20_f2_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f3_20_f3_20_f3_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f4_20_f4_20_f4_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f5_20_f5_20_f5_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f6_20_f6_20_f6_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f7_20_f7_20_f7_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f8_20_f8_20_f8_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_f9_20_f9_20_f9_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fa_20_fa_20_fa_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fb_20_fb_20_fb_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fc_20_fc_20_fc_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fd_20_fd_20_fd_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_fe_20_fe_20_fe_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		data_wen = 1'b1;
		//			   |<--				--->| |<--Ax---Ay----Az--T--->||<--Wx--Wy---Wz---T-->||<-Roll-Pit--Yaw--T-->|
		data_i = {256'h00_00_00_00_00_00_00_00_ff_20_ff_20_ff_20_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00, 1'b1};
		# 100;
		data_wen = 1'b0;
		# 39900;		// 400 - period
		end

	// ThresholdCutterWindow
	ThresholdCutterWindow #(
		.SIM_ENABLE(SIM_ENABLE),						// enable simulation
		.WINDOW_DEPTH_INDEX(WINDOW_DEPTH_INDEX),		// support up to 128 windows
		.WINDOW_DEPTH(WINDOW_DEPTH),					// 100 windows
		.WINDOW_WIDTH(WINDOW_WIDTH),					// 32-bit window
		.THRESHOLD(THRESHOLD),							// threshold
		.BLOCK_NUM_INDEX(BLOCK_NUM_INDEX),				// 2 ** 6 == 64 blocks
		.A_OFFSET(A_OFFSET),							// A's offset
		.SQUARE_SRC_DATA_WIDTH(SQUARE_SRC_DATA_WIDTH),	// square src data width
		.PRESET_SEQUENCE(PRESET_SEQUENCE)				// preset-sequence
	) m_ThresholdCutterWindow (
		.clk			(clk					),
		.rst_n			(rst_n					),

		.data_i			(data_i					),
		.data_wen		(data_wen				),

		.flag_o			(flag_o					)
	);

endmodule
