`timescale 1ns/1ns
module test_ThresholdCutterWindow #(
	`define			sim_window
) (

);

	

endmodule
