`timescale 1ns/1ns
module test_ThresholdCutter #(
	parameter		// config enable
					CONFIG_EN							=	0,		// do not enable config
					// config
					CLK_FRE								=	50,		// 50MHz
					BAUD_RATE							=	115200,	// 115200Hz (4800, 19200, 38400, 57600, 115200, 38400...)
					STOP_BIT							=	0,		// 0 : 1-bit stop-bit, 1 : 2-bit stop-bit
					CHECK_BIT							=	0,		// 0 : no check-bit, 1 : odd, 2 : even
					// default	9600	0	0
					// granularity
					REQUEST_FIFO_DATA_WIDTH				=	8,		// the bit width of data we stored in the FIFO
					REQUEST_FIFO_DATA_DEPTH_INDEX		=	6,		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
					RESPONSE_FIFO_DATA_WIDTH			=	8,		// the bit width of data we stored in the FIFO
					RESPONSE_FIFO_DATA_DEPTH_INDEX		=	6,		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
					// uart connected with PC
					PC_BAUD_RATE						=	115200,	// 115200Hz
					// enable simulation
					SIM_ENABLE							=	1,				// enable simulation
					// parameter for window
					WINDOW_DEPTH_INDEX					=	7,				// support up to 128 windows
					WINDOW_DEPTH						=	100,			// 100 windows
					WINDOW_WIDTH						=	(32 << 3),		// 32B window
					THRESHOLD							=	32'h0010_0000,	// threshold
					BLOCK_NUM_INDEX						=	4,				// 2 ** 6 == 64 blocks		// 16
					// parameter for package
					A_OFFSET							=	2,				// A's offset
					// parameter for square
					SQUARE_SRC_DATA_WIDTH				=	16,				// square src data width
					// parameter for preset-sequence
					PRESET_SEQUENCE						=	128'h00_01_02_03_04_05_06_07_08_09_00_01_02_03_04_05,
					// parameter for package
					PACKAGE_SIZE						=	11,
					PACKAGE_NUM							=	4,
					// parameter for uart
					TX_DATA_BYTE_WIDTH					=	11,		// 11 bytes to transmit
					RX_DATA_BYTE_WIDTH					=	11		// 11 bytes to receive
	`ifndef			TX_DATA_BIT_WIDTH
	`define			TX_DATA_BIT_WIDTH					(TX_DATA_BYTE_WIDTH << 3)
	`endif
	`ifndef			RX_DATA_BIT_WIDTH
	`define			RX_DATA_BIT_WIDTH					(RX_DATA_BYTE_WIDTH << 3)
	`endif
) (

);

	reg clk, rst_n;
	// ThresholdCutter signals
	wire BlueTooth_Txd;
	// sim_BlueTooth signals
	wire uart_tx;
	reg tx_vld;
	reg [`TX_DATA_BIT_WIDTH - 1:0] tx_data;

	// testsuite
	always # 50
		clk = ~clk;

	initial
		begin
		clk = 1'b0;
		rst_n = 1'b1;
		tx_vld = 1'b0;
		tx_data = {WINDOW_WIDTH{1'b0}};
		# 500;
		rst_n = 1'b0;
		# 500;
		rst_n = 1'b1;
		// begin
		/*
		tx_vld = 1'b1;
		tx_data = 88'h01_23_45_67_89_ab_cd_ef_fe_dc_ba;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h98_76_54_32_10_01_23_45_67_89_ab;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'hcd_ef_fe_dc_ba_98_76_54_32_10_01;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h23_45_67_89_ab_cd_ef_fe_dc_ba_98;
		*/
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_20_00_20_00_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_01_20_01_20_01_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_02_20_02_20_02_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_03_20_03_20_03_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_04_20_04_20_04_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_05_20_05_20_05_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_06_20_06_20_06_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_07_20_07_20_07_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_08_20_08_20_08_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_09_20_09_20_09_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0a_20_0a_20_0a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0b_20_0b_20_0b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0c_20_0c_20_0c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0d_20_0d_20_0d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0e_20_0e_20_0e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0f_20_0f_20_0f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_10_20_10_20_10_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_11_20_11_20_11_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_12_20_12_20_12_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_13_20_13_20_13_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_14_20_14_20_14_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_15_20_15_20_15_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_16_20_16_20_16_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_17_20_17_20_17_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_18_20_18_20_18_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_19_20_19_20_19_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1a_20_1a_20_1a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1b_20_1b_20_1b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1c_20_1c_20_1c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1d_20_1d_20_1d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1e_20_1e_20_1e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1f_20_1f_20_1f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_20_20_20_20_20_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_21_20_21_20_21_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_22_20_22_20_22_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_23_20_23_20_23_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_24_20_24_20_24_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_25_20_25_20_25_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_26_20_26_20_26_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_27_20_27_20_27_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_28_20_28_20_28_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_29_20_29_20_29_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2a_20_2a_20_2a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2b_20_2b_20_2b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2c_20_2c_20_2c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2d_20_2d_20_2d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2e_20_2e_20_2e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2f_20_2f_20_2f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_30_20_30_20_30_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_31_20_31_20_31_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_32_20_32_20_32_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_33_20_33_20_33_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_34_20_34_20_34_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_35_20_35_20_35_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_36_20_36_20_36_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_37_20_37_20_37_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_38_20_38_20_38_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_39_20_39_20_39_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3a_20_3a_20_3a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3b_20_3b_20_3b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3c_20_3c_20_3c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3d_20_3d_20_3d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3e_20_3e_20_3e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3f_20_3f_20_3f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_40_20_40_20_40_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_41_20_41_20_41_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_42_20_42_20_42_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_43_20_43_20_43_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_44_20_44_20_44_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_45_20_45_20_45_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_46_20_46_20_46_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_47_20_47_20_47_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_48_20_48_20_48_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_49_20_49_20_49_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4a_20_4a_20_4a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4b_20_4b_20_4b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4c_20_4c_20_4c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4d_20_4d_20_4d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4e_20_4e_20_4e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4f_20_4f_20_4f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_50_20_50_20_50_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_51_20_51_20_51_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_52_20_52_20_52_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_53_20_53_20_53_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_54_20_54_20_54_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_55_20_55_20_55_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_56_20_56_20_56_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_57_20_57_20_57_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_58_20_58_20_58_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_59_20_59_20_59_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5a_20_5a_20_5a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5b_20_5b_20_5b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5c_20_5c_20_5c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5d_20_5d_20_5d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5e_20_5e_20_5e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5f_20_5f_20_5f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_60_20_60_20_60_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_61_20_61_20_61_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_62_20_62_20_62_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_63_20_63_20_63_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_64_20_64_20_64_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_65_20_65_20_65_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_66_20_66_20_66_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_67_20_67_20_67_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_68_20_68_20_68_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_69_20_69_20_69_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6a_20_6a_20_6a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6b_20_6b_20_6b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6c_20_6c_20_6c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6d_20_6d_20_6d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6e_20_6e_20_6e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6f_20_6f_20_6f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_70_20_70_20_70_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_71_20_71_20_71_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_72_20_72_20_72_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_73_20_73_20_73_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_74_20_74_20_74_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_75_20_75_20_75_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_76_20_76_20_76_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_77_20_77_20_77_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_78_20_78_20_78_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_79_20_79_20_79_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7a_20_7a_20_7a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7b_20_7b_20_7b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7c_20_7c_20_7c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7d_20_7d_20_7d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7e_20_7e_20_7e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7f_20_7f_20_7f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_80_20_80_20_80_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_81_20_81_20_81_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_82_20_82_20_82_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_83_20_83_20_83_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_84_20_84_20_84_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_85_20_85_20_85_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_86_20_86_20_86_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_87_20_87_20_87_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_88_20_88_20_88_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_89_20_89_20_89_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8a_20_8a_20_8a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8b_20_8b_20_8b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8c_20_8c_20_8c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8d_20_8d_20_8d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8e_20_8e_20_8e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8f_20_8f_20_8f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_90_20_90_20_90_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_91_20_91_20_91_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_92_20_92_20_92_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_93_20_93_20_93_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_94_20_94_20_94_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_95_20_95_20_95_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_96_20_96_20_96_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_97_20_97_20_97_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_98_20_98_20_98_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_99_20_99_20_99_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9a_20_9a_20_9a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9b_20_9b_20_9b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9c_20_9c_20_9c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9d_20_9d_20_9d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9e_20_9e_20_9e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9f_20_9f_20_9f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a0_20_a0_20_a0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a1_20_a1_20_a1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a2_20_a2_20_a2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a3_20_a3_20_a3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a4_20_a4_20_a4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a5_20_a5_20_a5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a6_20_a6_20_a6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a7_20_a7_20_a7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a8_20_a8_20_a8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a9_20_a9_20_a9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_aa_20_aa_20_aa_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ab_20_ab_20_ab_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ac_20_ac_20_ac_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ad_20_ad_20_ad_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ae_20_ae_20_ae_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_af_20_af_20_af_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b0_20_b0_20_b0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b1_20_b1_20_b1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b2_20_b2_20_b2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b3_20_b3_20_b3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b4_20_b4_20_b4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b5_20_b5_20_b5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b6_20_b6_20_b6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b7_20_b7_20_b7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b8_20_b8_20_b8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b9_20_b9_20_b9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ba_20_ba_20_ba_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bb_20_bb_20_bb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bc_20_bc_20_bc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bd_20_bd_20_bd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_be_20_be_20_be_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bf_20_bf_20_bf_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c0_20_c0_20_c0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c1_20_c1_20_c1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c2_20_c2_20_c2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c3_20_c3_20_c3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c4_20_c4_20_c4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c5_20_c5_20_c5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c6_20_c6_20_c6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c7_20_c7_20_c7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c8_20_c8_20_c8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c9_20_c9_20_c9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ca_20_ca_20_ca_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cb_20_cb_20_cb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cc_20_cc_20_cc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cd_20_cd_20_cd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ce_20_ce_20_ce_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cf_20_cf_20_cf_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d0_20_d0_20_d0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d1_20_d1_20_d1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d2_20_d2_20_d2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d3_20_d3_20_d3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d4_20_d4_20_d4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d5_20_d5_20_d5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d6_20_d6_20_d6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d7_20_d7_20_d7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d8_20_d8_20_d8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d9_20_d9_20_d9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_da_20_da_20_da_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_db_20_db_20_db_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_dc_20_dc_20_dc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_dd_20_dd_20_dd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_de_20_de_20_de_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_df_20_df_20_df_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e0_20_e0_20_e0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e1_20_e1_20_e1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e2_20_e2_20_e2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e3_20_e3_20_e3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e4_20_e4_20_e4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e5_20_e5_20_e5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e6_20_e6_20_e6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e7_20_e7_20_e7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e8_20_e8_20_e8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e9_20_e9_20_e9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ea_20_ea_20_ea_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_eb_20_eb_20_eb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ec_20_ec_20_ec_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ed_20_ed_20_ed_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ee_20_ee_20_ee_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ef_20_ef_20_ef_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f0_20_f0_20_f0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f1_20_f1_20_f1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f2_20_f2_20_f2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f3_20_f3_20_f3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f4_20_f4_20_f4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f5_20_f5_20_f5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f6_20_f6_20_f6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f7_20_f7_20_f7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f8_20_f8_20_f8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f9_20_f9_20_f9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fa_20_fa_20_fa_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fb_20_fb_20_fb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fc_20_fc_20_fc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fd_20_fd_20_fd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fe_20_fe_20_fe_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ff_20_ff_20_ff_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_00_20_00_20_00_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_01_20_01_20_01_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_02_20_02_20_02_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_03_20_03_20_03_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_04_20_04_20_04_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_05_20_05_20_05_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_06_20_06_20_06_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_07_20_07_20_07_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_08_20_08_20_08_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_09_20_09_20_09_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0a_20_0a_20_0a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0b_20_0b_20_0b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0c_20_0c_20_0c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0d_20_0d_20_0d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0e_20_0e_20_0e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_0f_20_0f_20_0f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_10_20_10_20_10_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_11_20_11_20_11_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_12_20_12_20_12_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_13_20_13_20_13_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_14_20_14_20_14_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_15_20_15_20_15_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_16_20_16_20_16_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_17_20_17_20_17_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_18_20_18_20_18_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_19_20_19_20_19_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1a_20_1a_20_1a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1b_20_1b_20_1b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1c_20_1c_20_1c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1d_20_1d_20_1d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1e_20_1e_20_1e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_1f_20_1f_20_1f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_20_20_20_20_20_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_21_20_21_20_21_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_22_20_22_20_22_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_23_20_23_20_23_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_24_20_24_20_24_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_25_20_25_20_25_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_26_20_26_20_26_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_27_20_27_20_27_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_28_20_28_20_28_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_29_20_29_20_29_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2a_20_2a_20_2a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2b_20_2b_20_2b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2c_20_2c_20_2c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2d_20_2d_20_2d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2e_20_2e_20_2e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_2f_20_2f_20_2f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_30_20_30_20_30_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_31_20_31_20_31_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_32_20_32_20_32_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_33_20_33_20_33_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_34_20_34_20_34_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_35_20_35_20_35_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_36_20_36_20_36_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_37_20_37_20_37_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_38_20_38_20_38_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_39_20_39_20_39_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3a_20_3a_20_3a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3b_20_3b_20_3b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3c_20_3c_20_3c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3d_20_3d_20_3d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3e_20_3e_20_3e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_3f_20_3f_20_3f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_40_20_40_20_40_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_41_20_41_20_41_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_42_20_42_20_42_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_43_20_43_20_43_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_44_20_44_20_44_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_45_20_45_20_45_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_46_20_46_20_46_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_47_20_47_20_47_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_48_20_48_20_48_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_49_20_49_20_49_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4a_20_4a_20_4a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4b_20_4b_20_4b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4c_20_4c_20_4c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4d_20_4d_20_4d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4e_20_4e_20_4e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_4f_20_4f_20_4f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_50_20_50_20_50_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_51_20_51_20_51_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_52_20_52_20_52_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_53_20_53_20_53_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_54_20_54_20_54_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_55_20_55_20_55_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_56_20_56_20_56_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_57_20_57_20_57_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_58_20_58_20_58_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_59_20_59_20_59_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5a_20_5a_20_5a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5b_20_5b_20_5b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5c_20_5c_20_5c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5d_20_5d_20_5d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5e_20_5e_20_5e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_5f_20_5f_20_5f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_60_20_60_20_60_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_61_20_61_20_61_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_62_20_62_20_62_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_63_20_63_20_63_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_64_20_64_20_64_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_65_20_65_20_65_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_66_20_66_20_66_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_67_20_67_20_67_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_68_20_68_20_68_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_69_20_69_20_69_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6a_20_6a_20_6a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6b_20_6b_20_6b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6c_20_6c_20_6c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6d_20_6d_20_6d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6e_20_6e_20_6e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_6f_20_6f_20_6f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_70_20_70_20_70_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_71_20_71_20_71_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_72_20_72_20_72_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_73_20_73_20_73_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_74_20_74_20_74_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_75_20_75_20_75_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_76_20_76_20_76_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_77_20_77_20_77_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_78_20_78_20_78_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_79_20_79_20_79_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7a_20_7a_20_7a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7b_20_7b_20_7b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7c_20_7c_20_7c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7d_20_7d_20_7d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7e_20_7e_20_7e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_7f_20_7f_20_7f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_80_20_80_20_80_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_81_20_81_20_81_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_82_20_82_20_82_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_83_20_83_20_83_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_84_20_84_20_84_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_85_20_85_20_85_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_86_20_86_20_86_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_87_20_87_20_87_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_88_20_88_20_88_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_89_20_89_20_89_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8a_20_8a_20_8a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8b_20_8b_20_8b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8c_20_8c_20_8c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8d_20_8d_20_8d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8e_20_8e_20_8e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_8f_20_8f_20_8f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_90_20_90_20_90_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_91_20_91_20_91_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_92_20_92_20_92_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_93_20_93_20_93_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_94_20_94_20_94_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_95_20_95_20_95_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_96_20_96_20_96_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_97_20_97_20_97_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_98_20_98_20_98_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_99_20_99_20_99_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9a_20_9a_20_9a_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9b_20_9b_20_9b_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9c_20_9c_20_9c_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9d_20_9d_20_9d_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9e_20_9e_20_9e_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_9f_20_9f_20_9f_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a0_20_a0_20_a0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a1_20_a1_20_a1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a2_20_a2_20_a2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a3_20_a3_20_a3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a4_20_a4_20_a4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a5_20_a5_20_a5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a6_20_a6_20_a6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a7_20_a7_20_a7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a8_20_a8_20_a8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_a9_20_a9_20_a9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_aa_20_aa_20_aa_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ab_20_ab_20_ab_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ac_20_ac_20_ac_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ad_20_ad_20_ad_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ae_20_ae_20_ae_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_af_20_af_20_af_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b0_20_b0_20_b0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b1_20_b1_20_b1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b2_20_b2_20_b2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b3_20_b3_20_b3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b4_20_b4_20_b4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b5_20_b5_20_b5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b6_20_b6_20_b6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b7_20_b7_20_b7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b8_20_b8_20_b8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_b9_20_b9_20_b9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ba_20_ba_20_ba_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bb_20_bb_20_bb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bc_20_bc_20_bc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bd_20_bd_20_bd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_be_20_be_20_be_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_bf_20_bf_20_bf_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c0_20_c0_20_c0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c1_20_c1_20_c1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c2_20_c2_20_c2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c3_20_c3_20_c3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c4_20_c4_20_c4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c5_20_c5_20_c5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c6_20_c6_20_c6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c7_20_c7_20_c7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c8_20_c8_20_c8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_c9_20_c9_20_c9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ca_20_ca_20_ca_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cb_20_cb_20_cb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cc_20_cc_20_cc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cd_20_cd_20_cd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ce_20_ce_20_ce_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_cf_20_cf_20_cf_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d0_20_d0_20_d0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d1_20_d1_20_d1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d2_20_d2_20_d2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d3_20_d3_20_d3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d4_20_d4_20_d4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d5_20_d5_20_d5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d6_20_d6_20_d6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d7_20_d7_20_d7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d8_20_d8_20_d8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_d9_20_d9_20_d9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_da_20_da_20_da_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_db_20_db_20_db_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_dc_20_dc_20_dc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_dd_20_dd_20_dd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_de_20_de_20_de_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_df_20_df_20_df_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e0_20_e0_20_e0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e1_20_e1_20_e1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e2_20_e2_20_e2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e3_20_e3_20_e3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e4_20_e4_20_e4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e5_20_e5_20_e5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e6_20_e6_20_e6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e7_20_e7_20_e7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e8_20_e8_20_e8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_e9_20_e9_20_e9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ea_20_ea_20_ea_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_eb_20_eb_20_eb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ec_20_ec_20_ec_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ed_20_ed_20_ed_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ee_20_ee_20_ee_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ef_20_ef_20_ef_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f0_20_f0_20_f0_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f1_20_f1_20_f1_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f2_20_f2_20_f2_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f3_20_f3_20_f3_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f4_20_f4_20_f4_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f5_20_f5_20_f5_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f6_20_f6_20_f6_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f7_20_f7_20_f7_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f8_20_f8_20_f8_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_f9_20_f9_20_f9_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fa_20_fa_20_fa_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fb_20_fb_20_fb_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fc_20_fc_20_fc_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fd_20_fd_20_fd_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_fe_20_fe_20_fe_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_50_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_51_ff_20_ff_20_ff_20_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_52_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		tx_vld = 1'b1;
		tx_data = 88'h55_53_00_00_00_00_00_00_00_00_00;
		# 100;
		tx_vld = 1'b0;
		# 4999900;		// 400 - period
		end

	// sim_BlueTooth
	sim_BlueTooth #(
		// config
		.CLK_FRE(CLK_FRE),		// 50MHz
		.BAUD_RATE(BAUD_RATE),	// 9600Hz (4800, 19200, 38400, 57600, 115200, 38400...)
		.TX_DATA_BYTE_WIDTH(TX_DATA_BYTE_WIDTH),	// 11 bytes to transmit
		.RX_DATA_BYTE_WIDTH(RX_DATA_BYTE_WIDTH)		// 11 bytes to receive
	) m_sim_BlueTooth (
		.clk				(clk			),
		.rst_n				(rst_n			),

		// uart signals
		.uart_rx			(				),
		.uart_tx			(uart_tx		),		// should connect with BlueTooth_Txd in BlueToothController.v

		// inner data
		.tx_data			(tx_data		),		// data
		.tx_vld				(tx_vld			),		// start the transmit process
		.tx_rdy				(				),		// transmit process complete
		.rx_data			(				),		// data
		.rx_ack				(				),		// data is received by receiver buffer					(RX_WAIT)
		.rx_rdy				(				)		// send signal to receiver buffer that data is ready
	);

	// ThresholdCutter
	ThresholdCutter #(
		// config enable
		.CONFIG_EN(CONFIG_EN),		// do not enable config
		// config
		.CLK_FRE(CLK_FRE),		// 50MHz
		.BAUD_RATE(BAUD_RATE),	// 115200Hz (4800, 19200, 38400, 57600, 115200, 38400...)
		.STOP_BIT(STOP_BIT),		// 0 : 1-bit stop-bit, 1 : 2-bit stop-bit
		.CHECK_BIT(CHECK_BIT),		// 0 : no check-bit, 1 : odd, 2 : even
		// default	9600	0	0
		// granularity
		.REQUEST_FIFO_DATA_WIDTH(REQUEST_FIFO_DATA_WIDTH),		// the bit width of data we stored in the FIFO
		.REQUEST_FIFO_DATA_DEPTH_INDEX(REQUEST_FIFO_DATA_DEPTH_INDEX),		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
		.RESPONSE_FIFO_DATA_WIDTH(RESPONSE_FIFO_DATA_WIDTH),		// the bit width of data we stored in the FIFO
		.RESPONSE_FIFO_DATA_DEPTH_INDEX(RESPONSE_FIFO_DATA_DEPTH_INDEX),		// the index_width of data unit(reg [DATA_WIDTH - 1:0])
		// uart connected with PC
		.PC_BAUD_RATE(PC_BAUD_RATE),	// 115200Hz
		// enable simulation
		.SIM_ENABLE(SIM_ENABLE),				// enable simulation
		// parameter for window
		.WINDOW_DEPTH_INDEX(WINDOW_DEPTH_INDEX),				// support up to 128 windows
		.WINDOW_DEPTH(WINDOW_DEPTH),			// 100 windows
		.WINDOW_WIDTH(WINDOW_WIDTH),		// 32B window
		.THRESHOLD(THRESHOLD),	// threshold
		.BLOCK_NUM_INDEX(BLOCK_NUM_INDEX),				// 2 ** 6 == 64 blocks		// 16
		// parameter for package
		.A_OFFSET(A_OFFSET),				// A's offset
		// parameter for square
		.SQUARE_SRC_DATA_WIDTH(SQUARE_SRC_DATA_WIDTH),				// square src data width
		// parameter for preset-sequence
		.PRESET_SEQUENCE(PRESET_SEQUENCE),
		// parameter for package
		.PACKAGE_SIZE(PACKAGE_SIZE),
		.PACKAGE_NUM(PACKAGE_NUM)
	) m_ThresholdCutter (
		.clk							(clk				),
		.rst_n							(rst_n				),

		// BlueTooth_Config
		.BlueTooth_State				(					),
		.BlueTooth_Key					(					),
		.BlueTooth_Rxd					(					),
		.BlueTooth_Txd					(BlueTooth_Txd		),
		.BlueTooth_Vcc					(					),
		.BlueTooth_Gnd					(					),

		// ThresholdCutterWindow signals
		.ThresholdCutterWindow_flag_o	(					),

		// AXI RAM signals
		// ram safe access
		.rsta_busy						(					),
		.rstb_busy						(					),

		// AXI read control signals
		.s_axi_arid						(					),
		.s_axi_araddr					(					),
		.s_axi_arlen					(					),
		.s_axi_arsize					(					),
		.s_axi_arburst					(					),
		.s_axi_arvalid					(					),
		.s_axi_arready					(					),

		// AXI read data signals
		.s_axi_rid						(					),
		.s_axi_rdata					(					),
		.s_axi_rresp					(					),
		.s_axi_rlast					(					),
		.s_axi_rvalid					(					),
		.s_axi_rready					(					)
	);
	assign BlueTooth_Txd = uart_tx;

endmodule
